//-----------------------------------------------------------------------------
// 1-bit full_adde
//-----------------------------------------------------------------------------


module full_adder(in0, in1, cin, out, cout);
input in0, in1, cin;
output out, cout;

assign out = in0 ^ in1 ^ cin;
assign cout = ((in0 ^ in1) & cin) | (in0 & in1);
endmodule